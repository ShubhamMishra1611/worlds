module HelloWorld;
    initial begin
        $display("Hello, World!");
    end
endmodule